* SPICE3 file created from nandgate.ext - technology: scmos

.option scale=1u

M1000 vdd b z vdd pfet w=8 l=3
+  ad=168 pd=74 as=136 ps=50
M1001 z a vdd vdd pfet w=8 l=3
+  ad=0 pd=0 as=0 ps=0
M1002 z a gnd Gnd nfet w=8 l=3
+  ad=248 pd=94 as=56 ps=30
M1003 z b z Gnd nfet w=8 l=3
+  ad=0 pd=0 as=0 ps=0
C0 gnd Gnd 9.78fF
C1 z Gnd 6.39fF
C2 b Gnd 6.46fF
C3 a Gnd 6.46fF

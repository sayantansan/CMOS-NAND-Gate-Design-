magic
tech scmos
timestamp 1613423167
<< nwell >>
rect 0 0 46 25
<< polysilicon >>
rect 8 10 11 12
rect 28 10 31 12
rect 8 -3 11 2
rect 28 -1 31 2
rect 7 -7 11 -3
rect 27 -5 31 -1
rect 8 -13 11 -7
rect 28 -13 31 -5
rect 8 -23 11 -21
rect 28 -23 31 -21
<< ndiffusion >>
rect 1 -16 8 -13
rect 5 -20 8 -16
rect 1 -21 8 -20
rect 11 -15 28 -13
rect 11 -19 15 -15
rect 19 -19 28 -15
rect 11 -21 28 -19
rect 31 -14 45 -13
rect 31 -18 35 -14
rect 39 -18 45 -14
rect 31 -21 45 -18
<< pdiffusion >>
rect 5 6 8 10
rect 1 2 8 6
rect 11 8 28 10
rect 11 4 15 8
rect 19 4 28 8
rect 11 2 28 4
rect 31 6 34 10
rect 38 6 45 10
rect 31 2 45 6
<< metal1 >>
rect 4 16 9 20
rect 13 16 20 20
rect 24 16 31 20
rect 35 16 41 20
rect 45 16 46 20
rect 0 14 46 16
rect 1 10 5 14
rect 34 10 38 14
rect 15 8 19 9
rect 15 -8 19 4
rect 15 -12 44 -8
rect 15 -15 19 -12
rect 35 -14 39 -12
rect 1 -24 5 -20
rect 0 -26 46 -24
rect 0 -30 1 -26
rect 5 -30 12 -26
rect 16 -30 23 -26
rect 27 -30 33 -26
rect 37 -30 42 -26
<< ntransistor >>
rect 8 -21 11 -13
rect 28 -21 31 -13
<< ptransistor >>
rect 8 2 11 10
rect 28 2 31 10
<< polycontact >>
rect 3 -7 7 -3
rect 23 -5 27 -1
<< ndcontact >>
rect 1 -20 5 -16
rect 15 -19 19 -15
rect 35 -18 39 -14
<< pdcontact >>
rect 1 6 5 10
rect 15 4 19 8
rect 34 6 38 10
<< psubstratepcontact >>
rect 1 -30 5 -26
rect 12 -30 16 -26
rect 23 -30 27 -26
rect 33 -30 37 -26
rect 42 -30 46 -26
<< nsubstratencontact >>
rect 0 16 4 20
rect 9 16 13 20
rect 20 16 24 20
rect 31 16 35 20
rect 41 16 45 20
<< labels >>
rlabel metal1 16 16 16 16 1 vdd
rlabel polycontact 5 -5 5 -5 3 a
rlabel polycontact 25 -3 25 -3 1 b
rlabel metal1 42 -10 42 -10 7 z
rlabel metal1 19 -27 19 -27 1 gnd
<< end >>
